module testbench;
ClockGen cg (clock);
CPU c (clock);
endmodule 
